0
2 0 0 0 0 g 1 c 0 2 2 2 19 2
0 0 0 0 0 g c
0 0 0 0 0 g c
0 0 0 0 0 g c
1 3 5 7 4 5 0 2 5 7 0 8 0 10 5 7 1 11 4 8 1 3 5 7 3 3 0 2 1 2 1 8 3 10 1 9 3 9 
-1
