1
0 0 0 0 2 g c 1 1 9 1
0 0 0 0 1 g c 2 1 8 1
0 0 0 0 0 g c 3 1 7 1
0 0 0 0 1 g c 4 1 6 1
5 0 4 1 4 2 5 3 4 4 1 5 4 6 1 7 3 8 3 9 5 10 2 11 3 12 1 13 0 14 2 15 0 16 4 17 3 18 
-1
