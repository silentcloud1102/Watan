1
0 0 0 0 0 g c 20 1 22 1
0 0 0 0 0 g c 10 1 34 1
0 0 0 0 0 g c 13 1 0 1
0 0 0 0 0 g c 2 1 4 1
3 12 5 7 2 9 2 6 3 3 1 10 2 10 2 12 2 8 0 2 1 6 4 8 2 10 5 7 0 12 2 10 3 9 1 12 3 8 
-1
