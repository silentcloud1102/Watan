0
0 0 0 0 0 g c
0 0 0 0 0 g c
0 0 0 0 0 g c
0 0 0 0 0 g c
3 11 1 12 2 3 2 12 2 9 5 7 2 10 4 5 3 2 5 7 2 10 1 5 0 4 1 10 3 4 5 7 0 3 1 5 1 10 
-1
