4
1 2 1 1 1 g 4 12 c 18 3
0 1 0 1 1 g 7 13 19 c 6 1 25 2
2 4 0 0 2 g 1 8 c 30 1
2 1 0 1 0 g 9 c 14 1
0 3 1 10 4 5 1 4 5 7 3 10 0 10 4 12 0 3 4 8 0 6 1 8 3 3 4 11 1 2 4 6 3 10 2 9 0 12 
8
