3
0 0 0 0 0 g c 44 0 36 0
0 0 0 0 0 g c 50 0 24 0
0 0 0 0 0 g c 31 0 10 0
0 0 0 0 0 g c 13 0 8 0
3 5 1 11 3 5 2 10 3 4 0 12 2 11 3 2 0 9 0 6 3 3 4 4 3 11 2 6 1 3 1 2 0 8 1 9 1 5 
-1
